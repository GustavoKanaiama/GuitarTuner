`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 25.07.2025 17:32:45
// Design Name: 
// Module Name: twiddler_mod
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module twiddler_mod# (
parameter  WIDTH=16
)(
    input [WIDTH-1:0] k,
    input [WIDTH-1:0] n,
    
    output [WIDTH-1:0] twiddler_out_real,
    output [WIDTH-1:0] twiddler_out_imag
    );

real pi = 3.14;





    
    
    
endmodule
